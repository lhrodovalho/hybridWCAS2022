.subckt barth ip im op om vdd vss
  xap ip om vdd vss inv2_1
  xam im op vdd vss inv2_1
  xbp ip x  vdd vss inv1_1
  xbm im x  vdd vss inv1_1
  xc  x  x  vdd vss inv2_1
  xdp x  om vdd vss inv2_1
  xdm x  op vdd vss inv2_1
.ends

