* CMOS inverter-based single-ended amplifiers open-loop testbench

* Include SkyWater sky130 device models
.lib "/usr/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice" tt
.param mc_mm_switch=0

.include "../aux/array5v0.spice"
.include "../aux/inv.spice"
.include "nauta.spice"
.include "barth.spice"
.include "manf.spice"
.include "barthmanf.spice"
.include "barthnauta.spice"
.include "nautanauta.spice"
.include "nautavieru.spice"
.include "manfvieru.spice"

.param pVDD = 3.0
.param pC   = 10p

VDD  vdd 0 dc {pVDD}
VSS  vss 0 0
ECM  cm vss q vss 1
xa q q vdd vss inv2_4

vin in cm 0 ac 1

x0 xp0 xm0 op0 om0 vdd vss nauta
cxp0 in  xp0 1T
cxm0 in  xm0 1T
lop0 op0 xm0 1T
lom0 om0 xp0 1T
cop0 op0 cm  {pC}
com0 om0 cm  {pC}

x1 xp1 xm1 op1 om1 vdd vss barth
cxp1 in  xp1 1T
cxm1 in  xm1 1T
lop1 op1 xm1 1T
lom1 om1 xp1 1T
cop1 op1 cm  {pC}
com1 om1 cm  {pC}

x2 xp2 xm2 op2 om2 vdd vss manf
cxp2 in  xp2 1T
cxm2 in  xm2 1T
lop2 op2 xm2 1T
lom2 om2 xp2 1T
cop2 op2 cm  {pC}
com2 om2 cm  {pC}

x3 xm3 xp3 op3 om3 vdd vss barthnauta
cxp3 in  xp3 1T
cxm3 in  xm3 1T
lop3 op3 xm3 1T
lom3 om3 xp3 1T
cop3 op3 cm  {pC}
com3 om3 cm  {pC}

x4 xp4 xm4 op4 om4 vdd vss barthmanf
cxp4 in  xp4 1T
cxm4 in  xm4 1T
lop4 op4 xm4 1T
lom4 om4 xp4 1T
cop4 op4 cm  {pC}
com4 om4 cm  {pC}

x5 xp5 xm5 op5 om5 vdd vss nautanauta
cxp5 in  xp5 1T
cxm5 in  xm5 1T
lop5 op5 xm5 1T
lom5 om5 xp5 1T
cop5 op5 cm  {pC}
com5 om5 cm  {pC}

x6 xp6 xm6 op6 om6 vdd vss nautavieru
cxp6 in  xp6 1T
cxm6 in  xm6 1T
lop6 op6 xm6 1T
lom6 om6 xp6 1T
cop6 op6 cm  {pC}
com6 om6 cm  {pC}

x7 xp7 xm7 op7 om7 vdd vss manfvieru
cxp7 in  xp7 1T
cxm7 in  xm7 1T
lop7 op7 xm7 1T
lom7 om7 xp7 1T
cop7 op7 cm  {pC}
com7 om7 cm  {pC}

.option gmin=1e-15
.param dx = 1
.ac dec 100 1k 1T

.control
	run

	let av0 = dB((op0+om0)/2)
	let av1 = dB((op1+om1)/2)
	let av2 = dB((op2+om2)/2)
	let av3 = dB((op3+om3)/2)
	let av4 = dB((op4+om4)/2)
	let av5 = dB((op5+om5)/2)
	let av6 = dB((op6+om6)/2)
	let av7 = dB((op7+om7)/2)

	plot av0 av1 av2
	plot av0 av3 av4
	plot av5 av6 av7

	meas ac av0_1khz find av0 at=1k
	meas ac av1_1khz find av1 at=1k
	meas ac av2_1khz find av2 at=1k
	meas ac av3_1khz find av3 at=1k
	meas ac av4_1khz find av4 at=1k
	meas ac av5_1khz find av5 at=1k
	meas ac av6_1khz find av6 at=1k
	meas ac av7_1khz find av7 at=1k
	
	wrdata ../data/ac_cm_av.txt av0 av1 av2 av3 av4 av5 av6 av7
		
.endc

.end
